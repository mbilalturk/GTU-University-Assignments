library verilog;
use verilog.vl_types.all;
entity Tb is
end Tb;
